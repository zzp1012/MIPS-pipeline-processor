`timescale 1ns / 1ps

module instr_mem(instruction, read_addr);
    parameter word = 32;
    parameter byte = 8;
    parameter line = 42;
    
    input   [word - 1:0]    read_addr;
    output  [word - 1:0]    instruction;
    
    reg     [byte - 1:0]    mem[4*line - 1:0];
    reg     [word - 1:0]    instruction;
    integer                 n;
    
    initial begin
            for (n = 0; n < 4*line; n = n + 1) begin
                mem[n] = 0;
            end
            { mem[0], mem[1], mem[2], mem[3] } = 32'b00100000000010000000000000100000; // 1
            { mem[4], mem[5], mem[6], mem[7] } = 32'b00100000000010010000000000110111; // 2
            { mem[8], mem[9], mem[10], mem[11] } = 32'b00000001000010011000000000100100; // 3
            { mem[12], mem[13], mem[14], mem[15] } = 32'b00000001000010011000000000100101; // 4
            { mem[16], mem[17], mem[18], mem[19] } = 32'b10101100000100000000000000000100; // 5
            { mem[20], mem[21], mem[22], mem[23] } = 32'b10101100000010000000000000001000; // 6
            { mem[24], mem[25], mem[26], mem[27] } = 32'b00000001000010011000100000100000; // 7
            { mem[28], mem[29], mem[30], mem[31] } = 32'b00000001000010011001000000100010; // 8
            { mem[32], mem[33], mem[34], mem[35] } = 32'b00010010001100100000000000001001; // 9
            { mem[36], mem[37], mem[38], mem[39] } = 32'b10001100000100010000000000000100; // 10
            { mem[40], mem[41], mem[42], mem[43] } = 32'b10001100000100110000000000001000; // 13
            { mem[44], mem[45], mem[46], mem[47] } = 32'b00110010001100100000000001001000; // 11
            { mem[48], mem[49], mem[50], mem[51] } = 32'b00010010001100100000000000001001; // 12
            { mem[52], mem[53], mem[54], mem[55] } = 32'b00010010000100110000000000001010; // 14
            { mem[56], mem[57], mem[58], mem[59] } = 32'b00000010010100011010000000101010; // 15
            { mem[60], mem[61], mem[62], mem[63] } = 32'b00010010100000000000000000001111; // 16
            { mem[64], mem[65], mem[66], mem[67] } = 32'b00000010001000001001000000100000; // 17
            { mem[68], mem[69], mem[70], mem[71] } = 32'b00001000000000000000000000001110; // 18
            { mem[72], mem[73], mem[74], mem[75] } = 32'b00100000000010000000000000000000; // 19
            { mem[76], mem[77], mem[78], mem[79] } = 32'b00100000000010010000000000000000; // 20
            { mem[80], mem[81], mem[82], mem[83] } = 32'b00001000000000000000000000011111; // 21
            { mem[84], mem[85], mem[86], mem[87] } = 32'b00100000000010000000000000000001; // 22
            { mem[88], mem[89], mem[90], mem[91] } = 32'b00100000000010010000000000000001; // 23
            { mem[92], mem[93], mem[94], mem[95] } = 32'b00001000000000000000000000011111; // 24
            { mem[96], mem[97], mem[98], mem[99] } = 32'b00100000000010000000000000000010; // 25
            { mem[100], mem[101], mem[102], mem[103] } = 32'b00100000000010010000000000000010; // 26
            { mem[104], mem[105], mem[106], mem[107] } = 32'b00001000000000000000000000011111; // 27
            { mem[108], mem[109], mem[110], mem[111] } = 32'b00100000000010000000000000000011; // 28
            { mem[112], mem[113], mem[114], mem[115] } = 32'b00100000000010010000000000000011; // 29
            { mem[116], mem[117], mem[118], mem[119] } = 32'b00001000000000000000000000011111; // 30
            // $readmemb("D:/JI/2020 fall/VE370 Intro to Computer Organization/Projects/P2/InstructionMem_for_P2_Demo_bonus.txt", mem);
    end
    
    always @(read_addr) begin
        instruction = {mem[read_addr], mem[read_addr+1], mem[read_addr+2], mem[read_addr+3]};
    end
endmodule
